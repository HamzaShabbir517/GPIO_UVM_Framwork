// Declaration of GPIO defines

`define NUM_PINS 32
