// Declaration of Package
package gpio_test_lib_pkg;
	
	// Import UVM Package
	import uvm_pkg::*;
	
	// Include UVM Macros
	`include "uvm_macros.svh"
	
	// Import other packages
	// Import Envrionment 
	import gpio_apb_env_pkg::*;
	// Import Bus Agent
	import apb_agent_pkg::*;
	// Import Design
	import gpio_agent_pkg::*;
	// Import Register Model
	import gpio_apb_reg_pkg::*;
	// Import Bus Sequence 
	import gpio_bus_sequence_lib_pkg::*;
	// Import Virtual Sequence 
	import gpio_virtual_sequence_lib_pkg::*;
	
	
	// Include the test 
	`include "base_test.svh"
	`include "gpio_port_test.svh"
	`include "apb_test.svh"
	`include "gpio_reg_test.svh"
	`include "virtual_sequence_test.svh"
	
endpackage
