module hvl_top;

	// Import Packages
	import uvm_pkg::*;
	import gpio_test_lib_pkg::*;
	
	initial begin
		// RUN UVM Test
		run_test();
	end
	
endmodule

