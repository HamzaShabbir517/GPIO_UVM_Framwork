// Declaration of Package
package gpio_apb_env_pkg;

	// Import UVM Package
	import uvm_pkg::*;
	
	// Include UVM Macros
	`include "uvm_macros.svh"
	
	// Include other packages
	import apb_agent_pkg::*;
	import gpio_agent_pkg::*;
	import gpio_apb_reg_pkg::*;
	
	
	// Include GPIO Environment Config
	`include "gpio_apb_env_config.svh"
	
	// Include GPIO Environment
	`include "gpio_apb_environment.svh"
	
endpackage
