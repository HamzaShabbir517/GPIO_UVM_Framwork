// Declaration of AXI4 Lites defines

`define addr_width 32
`define data_width 32
