// Declaration of APB defines

`define PADDR_SIZE 32
`define PDATA_SIZE 32
